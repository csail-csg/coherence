
// Copyright (c) 2017 Massachusetts Institute of Technology
// 
// Permission is hereby granted, free of charge, to any person
// obtaining a copy of this software and associated documentation
// files (the "Software"), to deal in the Software without
// restriction, including without limitation the rights to use, copy,
// modify, merge, publish, distribute, sublicense, and/or sell copies
// of the Software, and to permit persons to whom the Software is
// furnished to do so, subject to the following conditions:
// 
// The above copyright notice and this permission notice shall be
// included in all copies or substantial portions of the Software.
// 
// THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND,
// EXPRESS OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
// MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND
// NONINFRINGEMENT. IN NO EVENT SHALL THE AUTHORS OR COPYRIGHT HOLDERS
// BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN
// ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN
// CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
// SOFTWARE.

import Types::*;
import CCTypes::*;
import FShow::*;

`ifdef CCSIZES_FILE
`include `CCSIZES_FILE
`else
staticAssert(False, "ERROR: CCSIZES_FILE undefined");
`endif

// Memory
//typedef 0 LgMemBankNum;
//typedef 1 MemChildNum; // number of child for each bank
//typedef Bit#(TLog#(MemChildNum)) MemChild;
//
//typedef 8 MemLdQSz;
//typedef 4 MemWrBSz;
//
//typedef Bit#(TLog#(DirCRqNum)) MemLdRqId; // XXX assume Mem connects to Dir

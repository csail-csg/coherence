// just to make things compile
`define rv64 True
`define m True
`define a True
`define f True
`define d True
`define sizeSup 1
`define NUM_CORES 1
`define NUM_EPOCHS 1
`define NUM_SPEC_TAGS 1
`define ROB_SIZE 1
`define LDQ_SIZE 1
`define STQ_SIZE 1
`define SB_SIZE 1
`define DRAMLLC_MAX_READS 1
`define LOG_BOOT_ROM_BYTES 12

// used for checking deadlock
`define LOG_DEADLOCK_CYCLES 26
